��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  Y9 jG     A3      �  9 *G     A2      �  �9 �G     A1      �  i9 zG     A0      �  YQ j_     B0      �  �Q �_     B1      �  	Q _     B2      �  IQ Z_     B3          0   0     ���  CLogicIn�� 	 CLatchKey  `a po          �� 	 CTerminal  xl y�                             td |l         ����     ��  pI �W          �  �T �i                             �L �T         ����     ��  �I �W          �  �T �i                             �L �T         ����     ��  �a �o          �  �l ��      
                       �d �l         ����     �� 	 CLogicOut�  ���                �            ��    "      ��     ��  ���       	        �            x�    $      ��     ��  ���      	 	        �            �     &      ��     ��  8�9       	        �            0@    (      ��     ��  x�y       	        �            p�    *      ��    ��  CXOR�  ����                �          �  p�q�                �          �  x�y�               �            l���    -      ��    +��  @�A�                �          �  0�1�                �          �  8�9�               �            ,�D�    1      ��    ��   I 0W       4   �  8T 9i                             4L <T     6    ����     ��  a  o       7   �  (l )�                             $d ,l     9    ����     ��  CAND�  L� a�                           �  L� a�                           �   � 5�                �            4� L�     <      ��    ��  `I pW       ?   �  xT yi                             tL |T     A    ����     ��  Pa `o       B   �  hl i�                             dd ll     D    ����     +��  x� y�                            �  h� i�                            �  pq               �            d� |    F      ��    ��  COR�   !               �          �  � !�                �          �  �� ��                �            ��     K      ��    :��  L0a1               �          �  L a!               �          �   (5)               �            4L4    O      ��    :��  h!i               �          �  X!Y               �          �  �`�a               �            �Tl    S      ��    I��  �8�9               �          �  �(�)               �          �  �0�1               �            �$�<    W      ��    +��  89%                           �  ()%                           �  0<1Q               �            $$<<    [      ��    :��  !	                          �  � !�                           �  � �               �            ��     _      ��    :��  T�i�                          �  T�i�                          �  (�=�               �            <�T�    c      ��    +��  ����                           �  x�y�                           �  ����               �            t���    g      ��    +��   ��                �          �  ����                �          �  ����     	          �            ���    k      ��    :��  ����               �          �  ����               �          �  ����               �            ����    o      ��    :��  �@�A     
                     �  �0�1                          �  �8�9               �            �,�D    s      ��    +��  �H�]                           �  �H�]      
                     �  �t��               �            �\�t    w      ��    I��  �p�q               �          �  �`�a               �          �  `hui               �            t\�t    {      ��        0   0     ���  CWire�� 
 CCrossOver  v�|�        h���      �  �h ��       �  x�y�       ���  v�|�        x� y�       �  �0�I       �  �h �1       �  �@�A     
 ���  �,�4        �� �A      
 ���  �,�4        �0�1      �  �� ��       �  �0�1      ���  n,t4        `0�1      �  �0��       ���  n,t4        p q�       �  @hA�       ���  .d4l         hAi      �  @hai      ���  .d4l        0X1�       ���  &� ,�          � 9�       �  8h 9�        �  ()       ���  &� ,�         (� )	       �  `� i�       ���  f� l�         h� i�        �  xh y�        ���  f� l�         `� y�       �  h� i�        �  x� y�        �   � !�        �  pq!       �  ` q!      �    !)       �  �8�a       �   X1Y      �  0P1Y       �  � �)       �  8� 9       �   )	      �  ����       �  h�y�      �   �)�      �   ��       �  ����      ���  ����        ���      ���  ����        ����       �  �@�I      
 �  �p��       �  �8�a           0   0     �    0   0         0   0       �   �   �   � " � " $ i $ & m & ( 3 ( * / * - � - . � . / / * 1 � 1 2 � 2 3 3 ( 6 6 � 9 9 � < < � = = � > � > A A � D D � F � F G � G H H � K K � L L � M � M O O � P P � Q � Q S S � T T � U � U W W � X X � Y � Y [ � [ \ � \ ] ] � _ _ � ` ` � a � a c c � d d � e � e g � g h � h i i $ k � k l � l m m & o o � p p � q � q s s � t t � u � u w � w x � x y y � { { � | | � } � } � � d �  � � h � �  � � w  � s � � �  � � � t � M " � Y � � O � � - � � � . � 1 � � S � � } � � � 2 � � ` � 6 � � \ � � 9 � < � � � D � A � � � = � � G � F > L H � P � K Q W U T � ] � a X � [ _ � � g c � � e � k p y � � o � � � � l � x { q u |            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V          ffffff�?      �? s 