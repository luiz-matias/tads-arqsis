��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  Y9 jG     A3      �  9 *G     A2      �  �9 �G     A1      �  i9 zG     A0      �  YQ j_     B0      �  �Q �_     B1      �  	Q _     B2      �  IQ Z_     B3          0   0     ���  CXOR�� 	 CTerminal  ����                           �  x�y�                           �  ����               �            t���          ��    �� 	 CLogicOut�  ���       	        �            x�          ��    ��  CLogicIn�� 	 CLatchKey  `a po          �  xl y�                             td |l         ����     ��  pI �W          �  �T �i                             �L �T     !    ����     ��  �I �W       "   �  �T �i                             �L �T     $    ����     ��  �a �o       %   �  �l ��      
                       �d �l     '    ����     ��  ���                �            ��    )      ��    ��  ���      	 	        �            �     +      ��    ��  8�9       	        �            0@    -      ��    ��  x�y       	        �            p�    /      ��    ��  ����                �          �  p�q�                �          �  x�y�               �            l���    1      ��    ��  @�A�                �          �  0�1�                �          �  8�9�               �            ,�D�    5      ��    ��   I 0W       8   �  8T 9i                             4L <T     :    ����     ��  a  o       ;   �  (l )�                             $d ,l     =    ����     ��  CAND�  L� a�                           �  L� a�                           �   � 5�                �            4� L�     @      ��    ��  `I pW       C   �  xT yi                             tL |T     E    ����     ��  Pa `o       F   �  hl i�                             dd ll     H    ����     ��  x� y�                            �  h� i�                            �  pq               �            d� |    J      ��    ��  COR�   !               �          �  � !�                �          �  �� ��                �            ��     O      ��    >��  L0a1               �          �  L a!               �          �   (5)               �            4L4    S      ��    >��  h!i               �          �  X!Y               �          �  �`�a               �            �Tl    W      ��    M��  �8�9               �          �  �(�)               �          �  �0�1               �            �$�<    [      ��    ��  89%                           �  ()%                           �  0<1Q               �            $$<<    _      ��    >��  !	                          �  � !�                           �  � �               �            ��     c      ��    >��  T�i�                          �  T�i�                          �  (�=�               �            <�T�    g      ��    ��   ��                �          �  ����                �          �  ����     	          �            ���    k      ��    >��  ����               �          �  ����               �          �  ����               �            ����    o      ��    >��  �@�A     
                     �  �0�1                          �  �8�9               �            �,�D    s      ��    ��  �H�]                           �  �H�]      
                     �  �t��               �            �\�t    w      ��    M��  �p�q               �          �  �`�a               �          �  `hui               �            t\�t    {      ��        0   0     ���  CWire  ����       �  x�y�       ��� 
 CCrossOver  v�|�        h���      �  �h ��       ���  v�|�        x� y�       �  �0�I       �  �h �1       �  �@�A     
 ���  �,�4        �� �A      
 ���  �,�4        �0�1      �  �� ��       �  �0�1      ���  n,t4        `0�1      �  �0��       ���  n,t4        p q�       �  @hA�       ���  .d4l         hAi      �  @hai      ���  .d4l        0X1�       ���  &� ,�          � 9�       �  8h 9�        �  ()       ���  &� ,�         (� )	       �  `� i�       ���  f� l�         h� i�        �  xh y�        ���  f� l�         `� y�       �  h� i�        �  x� y�        �   � !�        �  pq!       �  ` q!      �    !)       �  �8�a       �   X1Y      �  0P1Y       �  � �)       �  8� 9       �   )	      �  h�y�      �   �)�      �   ��       �  ����      ���  ����        ���      ���  ����        ����       �  �@�I      
 �  �p��       �  �8�a           0   0     �    0   0         0   0      �   �          � ! ! � $ $ � ' ' � ) � ) + m + - 7 - / 3 / 1 � 1 2 � 2 3 3 / 5 � 5 6 � 6 7 7 - : : � = = � @ @ � A A � B � B E E � H H � J � J K � K L L � O O � P P � Q � Q S S � T T � U � U W W � X X � Y � Y [ [ � \ \ � ] � ] _ � _ ` � ` a a � c c � d d � e � e g g � h h � i � i k � k l � l m m + o o � p p � q � q s s � t t � u � u w � w x � x y y � { { � | | � } � } �  �  � � h � ! � � �  � � w $ � s � � � ' � � � t � Q ) � ] � � S � � 1 � � � 2 � 5 � � W � � } � � � 6 � � d � : � � ` � � = � @ � � � H � E � � � A � � K � J B P L � T � O U [ Y X � a � e \ � _ c � g � � i � k p y � � o � � � � l � x { q u |            �$s�        @     +        @            @    "V  (      �P                
         $@      �? V               �? V         
         $@      �? V               �? V          ffffff�?      �? s 